----------------------------------------------------------------------------------
-- Company: 			ENSEIRB-Matmeca
-- Engineer:			Sylvain MARIEL & Thomas MOREAU
-- 
-- Create Date:		19:50:49 02/13/2013 
-- Design Name: 		Unit� de traitement
-- Module Name:		UniteTraitement - Behavioral 
-- Project Name: 		Processeur8bits
-- Target Devices:	Spartan 6
-- Tool versions: 
-- Description: 		Processeur 8 bits �l�mentaire � 4 instructions
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UAL is
end UAL;

architecture Behavioral of UAL is

begin


end Behavioral;

